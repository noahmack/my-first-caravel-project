magic
tech sky130A
magscale 1 2
timestamp 1729457247
<< locali >>
rect 728 1352 1506 1440
rect 728 1188 970 1352
rect 1482 1188 1506 1352
rect 728 1166 1506 1188
rect 728 1054 1512 1166
rect 734 480 906 1054
rect 1328 480 1512 1054
rect 734 444 1514 480
rect 736 196 1600 206
rect 732 182 1600 196
rect 732 -386 914 182
rect 1342 -386 1600 182
rect 732 -494 1600 -386
rect 732 -706 1002 -494
rect 1568 -706 1600 -494
rect 732 -784 1600 -706
<< viali >>
rect 970 1188 1482 1352
rect 1002 -706 1568 -494
<< metal1 >>
rect 728 1352 1508 1384
rect 728 1188 970 1352
rect 1482 1188 1508 1352
rect 728 1066 1508 1188
rect 978 762 1032 1066
rect 486 334 686 418
rect 1096 334 1126 936
rect 1190 788 1242 794
rect 1190 688 1258 788
rect 1206 354 1258 688
rect 1598 354 1798 430
rect 486 298 1146 334
rect 486 276 1148 298
rect 486 218 686 276
rect 1000 -202 1054 -54
rect 1000 -306 1048 -202
rect 1106 -266 1148 276
rect 1206 296 1798 354
rect 1206 -134 1258 296
rect 1598 230 1798 296
rect 1000 -380 1054 -306
rect 730 -494 1598 -380
rect 730 -706 1002 -494
rect 1568 -706 1598 -494
rect 730 -750 1598 -706
use sky130_fd_pr__nfet_g5v0d10v5_UNEQ2N  XM1
timestamp 1729455980
transform 1 0 1126 0 1 -98
box -278 -358 278 358
use sky130_fd_pr__pfet_g5v0d10v5_KLAZY6  XM3
timestamp 1729455980
transform 1 0 1112 0 1 767
box -308 -397 308 397
<< labels >>
flabel metal1 744 1180 944 1380 0 FreeSans 256 0 0 0 VDD
port 3 nsew
flabel metal1 770 -694 970 -494 0 FreeSans 256 0 0 0 VSS
port 2 nsew
flabel metal1 486 218 686 418 0 FreeSans 256 0 0 0 Vin
port 1 nsew
flabel metal1 1598 230 1798 430 0 FreeSans 256 0 0 0 Vout
port 0 nsew
<< end >>
