** sch_path: /home/noahmack/ChipISU/my-first-caravel-project/xschem/invTB.sch
**.subckt invTB
x1 VDD Vout Vin GND inverter
V1 Vin GND pulse(0 1.8 1ns 1ns 1ns 5ns 10ns)
V2 VDD GND 2.5
**** begin user architecture code

.param mc_mm_switch=0
.param mc_pr_switch=0
.include /home/noahmack/ChipISU/my-first-caravel-project/dependencies/pdks/sky130A/libs.tech/ngspice/corners/tt.spice
.include /home/noahmack/ChipISU/my-first-caravel-project/dependencies/pdks/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical.spice
.include /home/noahmack/ChipISU/my-first-caravel-project/dependencies/pdks/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical__lin.spice
.include /home/noahmack/ChipISU/my-first-caravel-project/dependencies/pdks/sky130A/libs.tech/ngspice/corners/tt/specialized_cells.spice


.tran .01n 1u
.save all

**** end user architecture code
**.ends

* expanding   symbol:  inverter.sym # of pins=4
** sym_path: /home/noahmack/ChipISU/my-first-caravel-project/xschem/inverter.sym
** sch_path: /home/noahmack/ChipISU/my-first-caravel-project/xschem/inverter.sch
.subckt inverter VDD Vout Vin VSS
*.opin Vout
*.ipin Vin
*.iopin VSS
*.iopin VDD
XM3 Vout Vin VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM1 Vout Vin VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends

.GLOBAL GND
.end
