** sch_path: /home/noahmack/ChipISU/my-first-caravel-project/xschem/inverter.sch
.subckt inverter Vout Vin VSS VDD
*.PININFO Vout:O Vin:I VSS:B VDD:B
XM3 Vout Vin VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=1 nf=1 m=1
XM1 Vout Vin VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 m=1
.ends
.end
