* NGSPICE file created from inverter_flat.ext - technology: sky130A

.subckt inverter_flat Vout Vin VSS VDD
X0 Vout.t0 Vin.t0 VDD.t1 VDD.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1 Vout.t1 Vin.t1 VSS.t1 VSS.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
R0 Vin.n0 Vin.t0 121.54
R1 Vin.n0 Vin.t1 118.879
R2 Vin Vin.n0 1.04145
R3 VDD.n8 VDD.n7 955.241
R4 VDD.n5 VDD.n3 955.241
R5 VDD.n11 VDD.t1 227.966
R6 VDD.n3 VDD.n2 209.46
R7 VDD.n7 VDD.n6 209.46
R8 VDD.n4 VDD.n1 87.4018
R9 VDD.n4 VDD.n0 85.6441
R10 VDD.n5 VDD.n4 46.2505
R11 VDD.n9 VDD.n8 46.2505
R12 VDD.n8 VDD.n2 34.4421
R13 VDD.n6 VDD.n5 34.4421
R14 VDD.n9 VDD.n1 29.5125
R15 VDD.n3 VDD.n0 26.4581
R16 VDD.n7 VDD.n1 26.4291
R17 VDD.n10 VDD.n0 23.9398
R18 VDD.n6 VDD.t0 10.1424
R19 VDD.t0 VDD.n2 10.1424
R20 VDD.n10 VDD.n9 3.76132
R21 VDD.n11 VDD.n10 0.751657
R22 VDD VDD.n11 0.103094
R23 Vout.n0 Vout.t0 228.237
R24 Vout.n0 Vout.t1 83.7184
R25 Vout Vout.n0 0.848668
R26 VSS.n6 VSS.n2 1570.81
R27 VSS.n6 VSS.n3 1570.81
R28 VSS.n7 VSS.n3 1570.81
R29 VSS.n7 VSS.n2 1570.81
R30 VSS.n4 VSS.n2 874.211
R31 VSS.n4 VSS.n3 874.211
R32 VSS.n6 VSS.n5 146.25
R33 VSS.t0 VSS.n6 146.25
R34 VSS.n8 VSS.n7 146.25
R35 VSS.n7 VSS.t0 146.25
R36 VSS.n2 VSS.n0 97.5005
R37 VSS.n3 VSS.n1 97.5005
R38 VSS.n5 VSS.n1 92.213
R39 VSS.n5 VSS.n0 87.1412
R40 VSS.n10 VSS.t1 83.4771
R41 VSS.n8 VSS.n1 27.0527
R42 VSS.n9 VSS.n0 18.203
R43 VSS.t0 VSS.n4 17.7119
R44 VSS.n9 VSS.n8 4.9644
R45 VSS.n10 VSS.n9 0.475162
R46 VSS VSS.n10 0.0873243
C0 Vin VDD 0.596579f
C1 Vout Vin 0.486458f
C2 Vout VDD 0.285893f
C3 Vout VSS 0.62354f
C4 Vin VSS 1.07368f
C5 VDD VSS 2.84012f
.ends

